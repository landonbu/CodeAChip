module MovementDetect(one,two);
	input one;
	output two;
	assign two = one;
endmodule 